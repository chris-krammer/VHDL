--------------------------------------------------------------------------------------------------
--																								--
-- 																								--
-- 				F A C H H O C H S C H U L E 	- 	T E C H N I K U M W I E N					--
-- 																								--
-- 						 																		--
--------------------------------------------------------------------------------------------------
--																								--
-- Web: http://www.technikum-wien.at/															--
-- 																								--
-- Contact: christopher.krammer@technikum-wien.at												--
--																								--
--------------------------------------------------------------------------------------------------
--
--
-- Author: Christopher Krammer
--
-- Filename: counter_.vhd
--
-- Date of Creation: Sun Dec 16 21:33:00 2018
--
-- Version: 1.0
--
-- Date of Latest Version: Sun Dec 16 21:33:00 2018
--
-- Design Unit: counter (Configuration)
--
-- Description: Counts either up or down.
--				Min and Max values can be changed by generics.
--				Max Countvalue is restricted to 
--
--		!! Keep in Mind: Counting is NOT triggered by CLK_i (MasterClock)	!!		
--		!! Keep in Mind: Counting is triggered by SCLK_i (SlowClock)		!!
--
--------------------------------------------------------------------------------------------------
--
-- CVS Change Log:
--
--
--------------------------------------------------------------------------------------------------
configuration counter_fsm_rtl_cfg of counter_fsm is
  for rtl        -- architecture rtl is used for entity orgate
  end for;
end counter_fsm_rtl_cfg;