--------------------------------------------------------------------------------------------------
--                                                                                              --
--                                                                                              --
--                  F A C H H O C H S C H U L E   -   T E C H N I K U M W I E N                 --
--                                                                                              --
--                                                                                              --
--------------------------------------------------------------------------------------------------
--                                                                                              --
-- Web: http://www.technikum-wien.at/                                                           --
--                                                                                              --
-- Contact: es19m001@technikum-wien.at                                                          --
--------------------------------------------------------------------------------------------------
-- Author: Christopher Krammer
--
-- Filename: uart_rtl_cfg.vhd
--
-- Date of Creation: Wed Sep 04 07:30:00 2019
--
-- Version: 1.0
--
-- Date of Creation: Wed Sep 04 07:30:00 2019
--
-- Design Unit: uart (Configuration)
--
-- Description: UART Entity for Asynchronous communication
--------------------------------------------------------------------------------------------------
-- CVS Change Log:
--
--------------------------------------------------------------------------------------------------
configuration uart_rtl_cfg of uart is
  for rtl        -- architecture rtl is used for entity
  end for;
end uart_rtl_cfg;
