--------------------------------------------------------------------------------
--                                                                            --
--        F A C H H O C H S C H U L E   -   T E C H N I K U M W I E N         --
--                                                                            --
--------------------------------------------------------------------------------
--                                                                            --
-- Web: http://www.technikum-wien.at/                                         --
--                                                                            --
-- Contact: christopher.krammer@technikum-wien.at                             --
--                                                                            --
--------------------------------------------------------------------------------
--
-- Author: Christopher Krammer
--
-- Filename: mux4to1_rtl_cfg.vhd
--
-- Version: 1.0
--
-- Design Unit: mux4to1 (Configuration)
--
-- Description: Selects one of the four inputs and copies it to the output
--
--------------------------------------------------------------------------------
-- CVS Change Log:
--
--------------------------------------------------------------------------------
configuration mux4to1_rtl_cfg of mux4to1 is
  for rtl        -- architecture rtl is used for entity orgate
  end for;
end mux4to1_rtl_cfg;