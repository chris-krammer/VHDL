--------------------------------------------------------------------------------------------------
--                                                                                              --
--                                                                                              --
--                  F A C H H O C H S C H U L E   -   T E C H N I K U M W I E N                 --
--                                                                                              --
--                                                                                              --
--------------------------------------------------------------------------------------------------
--                                                                                              --
-- Web: http://www.technikum-wien.at/                                                           --
--                                                                                              --
-- Contact: christopher.krammer@technikum-wien.at                                               --
--------------------------------------------------------------------------------------------------
--
--
-- Author: Christopher Krammer
--
-- Filename: ioCtrl_rtl.vhd
--
-- Date of Creation: Sun Dec 16 21:33:00 2018
--
-- Version: 1.0
--
-- Date of Latest Version: Sun Dec 16 21:33:00 2018
--
-- Design Unit: mux4to1 (Architecture)
--
-- Description: Syncs and debounces the inputs and acts as last instance before outputs interact
--              with the "real" world
--------------------------------------------------------------------------------------------------
--
-- CVS Change Log:
--
--
--------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

architecture rtl of ioCtrl is
  -- Signals for 7-Segment Display
  signal s_SS_CLK_EN  : std_logic := '0';
  signal s_sel        : std_logic_vector( 1 downto 0) := (others => '0');
  signal s_ss_sel     : std_logic_vector( 3 downto 0) := (others => '0');
  signal s_ss         : std_logic_vector( 7 downto 0) := (others => '0');

  -- Used to generate 4 kHz clock for 7-Segment
  component clkPrescale is
    generic(g_SOURCEHZ  : integer   := 100e6;  -- Frequency of the Master Clock HZ
            g_TARGETHZ  : integer   :=   1e3;  -- Desired Frequency in HZ
            g_OUTACTIVE : std_logic :=   '1';  -- Defines ACTIVE state of output
            g_RSTACTIVE : std_logic :=   '0'   -- Defines ACTIVE state for RST_i
          );
    port(
      -- Inputs
      CLK_i : in std_logic;
      RST_i : in std_logic;
      -- Outputs
      OUT_o: out std_logic
      );
  end component clkPrescale;

  -- Used to mux through the 7-Segment digits and values
  component mux4to1 is
    generic(DataWidth : integer);  -- Define DataWidth of Input- and Output Signals
    port (
    -- Inputs
    IN0_i : in std_logic_vector(DataWidth - 1 downto 0);  -- Input 1
    IN1_i : in std_logic_vector(DataWidth - 1 downto 0);  -- Input 2
    IN2_i : in std_logic_vector(DataWidth - 1 downto 0);  -- Input 3
    IN3_i : in std_logic_vector(DataWidth - 1 downto 0);  -- Input 4
    SEL_i : in std_logic_vector(1 downto 0);  -- Input Select Signal
    -- Outputs
    OUT_o : out std_logic_vector(DataWidth - 1 downto 0)  -- Output
  );
  end component mux4to1;

  -- Used to debounce pushbuttons and switches for further internal use
  component debouncer is
    generic(  g_SOURCEHZ      : integer range 1 to 100e6 := 100e6;  -- Board Clock Frequency in Hz
              g_DEBTIME       : integer range 1 to 100 := 10;       -- Debounce Time in ms
              g_RSTACTIVE     : std_logic := '1'                    -- Reset ACTIVE state
            );
    port(
          --  Inputs
          CLK_i : in std_logic;  -- Board Clock
          RST_i : in std_logic;  -- Reset
          IN_i  : in std_logic;  -- Input to be debounced
          -- Outputs
          OUT_o : out std_logic
        );
  end component debouncer;

  ---------------------------------------------------------------------------------
  -- Function to set the correct segments based on the ioCtrl value
  ---------------------------------------------------------------------------------
  function SS_Val(CalcVal : std_logic_vector(3 downto 0)) return std_logic_vector is
  begin
  case CalcVal is
    when x"0" =>  return b"00000011";
    when x"1" =>  return b"10011111";
    when x"2" =>  return b"00100101";
    when x"3" =>  return b"00001101";
    when x"4" =>  return b"10011001";
    when x"5" =>  return b"01001001";
    when x"6" =>  return b"01000001";
    when x"7" =>  return b"00011111";
    when x"8" =>  return b"00000001";
    when x"9" =>  return b"00001001";
    when x"A" =>  return b"00010001";
    when x"B" =>  return b"11000001";
    when x"C" =>  return b"01100011";
    when x"D" =>  return b"10000101";
    when x"E" =>  return b"01100001";
    when x"F" =>  return b"01110001";
    when others => return x"FF"; -- All OFF
    end case;
  end function SS_Val;


begin -- rtl
  -----------------------------------------------------------------------------
  -- Debounce buttons and switches
  -- Debounces each element of the vector on its own
  -----------------------------------------------------------------------------
    GEN_PB_DEBOUNCER : for i in 0 to (g_PBINPUTS - 1) generate
      --PB_DEBx : entity work.debouncer(rtl)
      PB_DEBx : debouncer
        generic map(
          g_SOURCEHZ  => g_SOURCEHZ,
          g_DEBTIME   => g_DEBTIME,
          g_RSTACTIVE => g_RSTACTIVE
          )
        port map(
          CLK_i => CLK_i,
          RST_i => RST_i,
          IN_i  => PB_i(i),
          OUT_o => PBSYNC_o(i)
          );
    end generate GEN_PB_DEBOUNCER;

    GEN_SW_DEBOUNCER : for i in 0 to (g_SWINPUTS - 1) generate
      --SW_DEBx : entity work.debouncer(rtl)
      SW_DEBx : debouncer
        generic map(
          g_SOURCEHZ  => g_SOURCEHZ,
          g_DEBTIME   => g_DEBTIME,
          g_RSTACTIVE => g_RSTACTIVE
          )
        port map(
          CLK_i => CLK_i,
          RST_i => RST_i,
          IN_i  => SW_i(i),
          OUT_o => SWSYNC_o(i)
          );
    end generate GEN_SW_DEBOUNCER;

  ----------------------------------------------------------------------------
  -- Display controller for the 7-segment display
  -- Segment is ACTIVE when Signal is LOW!!
  -----------------------------------------------------------------------------
    -----------------------------------------------------------------------------
    -- 7-Segment Clock
    --   Fastest Counting Freq = 1 kHz = Period of 7-Segment
    --   -> each of the 4 7-Segments should be lit once per Period
    --   -> 4 * 1 kHz => 4 kHz Clock needed
    -----------------------------------------------------------------------------
    SS_Clock : clkPrescale
      generic map(  g_SOURCEHZ  =>  g_SOURCEHZ,
                    g_TARGETHZ  =>  4 * 1e3, -- 4kHz
                    g_OUTACTIVE =>  '1',
                    g_RSTACTIVE =>  g_RSTACTIVE
                  )

      port map( CLK_i => CLK_i,
                RST_i => RST_i,
                OUT_o => s_SS_CLK_EN
              );
    -----------------------------------------------------------------------------
    -- SELECT Generator for MUX (2 bit select)
    -- 00 -> 01 -> 10 -> 11 -> 00 ..
    -----------------------------------------------------------------------------
    p_displaycontrol : process (CLK_i)
    begin -- process displaycontroler

      -- Reset condition is not needed here,
      -- since during the RESET segments need to display 'nothing' (b"11111111")

      if (rising_edge(CLK_i)) then -- rising clock edge
        if s_SS_CLK_EN = '1' then
          s_sel <= std_logic_vector(unsigned(s_sel) + 1 );
        end if;
      end if;

    end process p_displaycontrol;

    -----------------------------------------------------------------------------
    -- DIGIT VALUE MUX - Controlled by p_displaycontrol
    -- Fetches the correct translation depending on the input signal
    -----------------------------------------------------------------------------
    SS_VALUE_SEL : mux4to1
      generic map (DataWidth => 8)
      port map( IN0_i => SS_Val(CNTR0_i),
                IN1_i => SS_Val(CNTR1_i),
                IN2_i => SS_Val(CNTR2_i),
                IN3_i => SS_Val(CNTR3_i),
                SEL_i => s_sel,
                OUT_o => s_ss
              );

    -----------------------------------------------------------------------------
    -- DIGIT SEL MUX - Controlled by p_displaycontrol
    -- Enables the corresponding digit on the 7-Segment
    -----------------------------------------------------------------------------
    SS_DIGIT_SEL : mux4to1
      generic map (DataWidth => 4)
      port map( IN0_i => b"1110",
                IN1_i => b"1101",
                IN2_i => b"1011",
                IN3_i => b"0111",
                SEL_i => s_sel,
                OUT_o => s_ss_sel
              );

    SS_o <= s_ss when RST_i = '0' else x"FF";
    SS_SEL_o <= s_ss_sel; -- Keep muxing even when reseted
  ----------------------------------------------------------------------------


end rtl;
